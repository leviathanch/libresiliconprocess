* Qucs 0.0.20 /home/leviathan/libresiliconprocess/simulation/1xinv.sch
.INCLUDE "/usr/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 0.0.20  /home/leviathan/libresiliconprocess/simulation/1xinv.sch
.INCLUDE "/home/leviathan/libresiliconprocess/simulation/pmos1u.lib"
.INCLUDE "/home/leviathan/libresiliconprocess/simulation/nmos1u.lib"
V3 _net0 0 DC 5
V2 _net1 0 DC 0 PULSE( 0  5 0N 100N 100N 1e-06 2.2e-06)  AC 0
EPr1 Pr1 0 output 0 1.0
XPMOS  output input _net0 _net0 LV1UPMOS 
R4 input _net1  50
R5 0 output  100K
XNMOS  output input 0 0 LV1UNMOS 
.control
echo "" > spice4qucs.cir.noise
echo "" > spice4qucs.cir.pz
tran 5e-08 1e-05 0 
write 1xinv_tran.txt v(Pr1) v(input) v(output) 
destroy all
reset

exit
.endc
.END
