magic
tech ls1u
timestamp 1531674388
<< nwell >>
rect 0 32 16 48
<< end >>
