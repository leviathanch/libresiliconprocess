magic
magscale 1 2
timestamp 1522775789716
<< pads >>
rect 1 1 181 181
rect 1 265 181 445
<< end >>
