magic
magscale 1 2
timestamp 1522784296024
<< poly >>
rect 1 1 181 181 
<< end >>
